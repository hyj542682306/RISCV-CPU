`include "Definition.v"

module Mem_ctrl (
	
);

endmodule //Mem_ctrl